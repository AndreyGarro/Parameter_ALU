module display #(parameter n=8) (input logic [n-1:0] in_hex,
											output logic [7:0] disp);
											
	
	
endmodule
