module test();

	logic [3:0] a, b; 
	logic [3:0] s;
	logic [3:0] c;
	logic zero, negative, _carry, overflow;

	param_alu #(4) DUT(a,b,s,c,zero, negative, _carry, overflow);

	initial begin
		s = 4'b0000;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b0001;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b0010;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b0011;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b0100;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b0101;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b1000;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b1001;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b1010;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
		
		#10 s = 4'b1011;
		a = 4'b1100; b = 4'b1010; 
		#10 a = 4'b1100; b = 4'b1010;
		#10 a = 4'b1101; b = 4'b1011;
	end
	
endmodule
